module coreir_ult #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 < in1;

endmodule  // coreir_ult

module coreir_reg #(parameter clk_posedge=1, parameter init=1, parameter width=1) (
  input clk,
  input [width-1:0] in,
  output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;

endmodule  // coreir_reg

module coreir_mux #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  input sel,
  output [width-1:0] out
);
  assign out = sel ? in1 : in0;

endmodule  // coreir_mux

module coreir_mul #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 * in1;

endmodule  // coreir_mul

module coreir_mem #(parameter depth=1, parameter has_init=0, parameter width=1) (
  input clk,
  input [width-1:0] wdata,
  input [$clog2(depth)-1:0] waddr,
  input wen,
  output [width-1:0] rdata,
  input [$clog2(depth)-1:0] raddr
);
  reg [width-1:0] data[depth-1:0];
  always @(posedge clk) begin
    if (wen) begin
      data[waddr] <= wdata;
    end
  end
  assign rdata = data[raddr];

endmodule  // coreir_mem

module coreir_eq #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 == in1;

endmodule  // coreir_eq

module coreir_const #(parameter value=1, parameter width=1) (
  output [width-1:0] out
);
  assign out = value;

endmodule  // coreir_const

module coreir_add #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 + in1;

endmodule  // coreir_add

module corebit_const #(parameter value=1) (
  output out
);
  assign out = value;

endmodule  // corebit_const

module corebit_and (
  input in0,
  input in1,
  output out
);
  assign out = in0 & in1;

endmodule  // corebit_and

module partialParallel2Convolution_Circuit (
  input  CE,
  input  CLK,
  input [7:0] I0,
  input [7:0] I1,
  output [7:0] O0,
  output [7:0] O1,
  output  ready_data_in,
  input  ready_data_out,
  input  valid_data_in,
  output  valid_data_out
);


  // Instancing generated Module: coreir.add(width:8)
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_0_0$coreir_add8_inst0__in0;
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_0_0$coreir_add8_inst0__in1;
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_0_0$coreir_add8_inst0__out;
  coreir_add #(.width(8)) ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_0_0$coreir_add8_inst0(
    .in0(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_0_0$coreir_add8_inst0__in0),
    .in1(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_0_0$coreir_add8_inst0__in1),
    .out(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_0_0$coreir_add8_inst0__out)
  );

  // Instancing generated Module: coreir.add(width:8)
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_0$coreir_add8_inst0__in0;
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_0$coreir_add8_inst0__in1;
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_0$coreir_add8_inst0__out;
  coreir_add #(.width(8)) ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_0$coreir_add8_inst0(
    .in0(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_0$coreir_add8_inst0__in0),
    .in1(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_0$coreir_add8_inst0__in1),
    .out(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_0$coreir_add8_inst0__out)
  );

  // Instancing generated Module: coreir.add(width:8)
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_1$coreir_add8_inst0__in0;
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_1$coreir_add8_inst0__in1;
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_1$coreir_add8_inst0__out;
  coreir_add #(.width(8)) ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_1$coreir_add8_inst0(
    .in0(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_1$coreir_add8_inst0__in0),
    .in1(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_1$coreir_add8_inst0__in1),
    .out(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_1$coreir_add8_inst0__out)
  );

  // Instancing generated Module: coreir.add(width:8)
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_0_0$coreir_add8_inst0__in0;
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_0_0$coreir_add8_inst0__in1;
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_0_0$coreir_add8_inst0__out;
  coreir_add #(.width(8)) ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_0_0$coreir_add8_inst0(
    .in0(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_0_0$coreir_add8_inst0__in0),
    .in1(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_0_0$coreir_add8_inst0__in1),
    .out(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_0_0$coreir_add8_inst0__out)
  );

  // Instancing generated Module: coreir.add(width:8)
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_0$coreir_add8_inst0__in0;
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_0$coreir_add8_inst0__in1;
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_0$coreir_add8_inst0__out;
  coreir_add #(.width(8)) ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_0$coreir_add8_inst0(
    .in0(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_0$coreir_add8_inst0__in0),
    .in1(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_0$coreir_add8_inst0__in1),
    .out(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_0$coreir_add8_inst0__out)
  );

  // Instancing generated Module: coreir.add(width:8)
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_1$coreir_add8_inst0__in0;
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_1$coreir_add8_inst0__in1;
  wire [7:0] ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_1$coreir_add8_inst0__out;
  coreir_add #(.width(8)) ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_1$coreir_add8_inst0(
    .in0(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_1$coreir_add8_inst0__in0),
    .in1(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_1$coreir_add8_inst0__in1),
    .out(ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_1$coreir_add8_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:3)
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join__in0;
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join__in1;
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join__sel;
  coreir_mux #(.width(3)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.const(width:3)
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$const_0_3__out;
  coreir_const #(.value(3'h0),.width(3)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$const_0_3(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$const_0_3__out)
  );

  // Instancing generated Module: coreir.mux(width:3)
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join__in0;
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join__in1;
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join__sel;
  coreir_mux #(.width(3)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:3)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__clk;
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__in;
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__out;
  coreir_reg #(.clk_posedge(1),.init(3'h0),.width(3)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__out)
  );

  // Instancing generated Module: coreir.const(width:3)
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$const_1_3__out;
  coreir_const #(.value(3'h1),.width(3)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$const_1_3(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$const_1_3__out)
  );

  // Instancing generated Module: coreir.add(width:3)
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$coreir_add3_inst0__in0;
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$coreir_add3_inst0__in1;
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$coreir_add3_inst0__out;
  coreir_add #(.width(3)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$coreir_add3_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$coreir_add3_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$coreir_add3_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$coreir_add3_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$and_inst0__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$and_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$and_inst0__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$and_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$and_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$and_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:3)
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$const_6_3__out;
  coreir_const #(.value(3'h6),.width(3)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$const_6_3(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$const_6_3__out)
  );

  // Instancing generated Module: coreir.eq(width:3)
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$coreir_eq_3_inst0__in0;
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$coreir_eq_3_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$coreir_eq_3_inst0__out;
  coreir_eq #(.width(3)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$coreir_eq_3_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$coreir_eq_3_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$coreir_eq_3_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$coreir_eq_3_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1__out;
  coreir_const #(.value(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$const_1_1__out;
  coreir_const #(.value(1'h1),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$const_1_1(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$const_1_1__out)
  );

  // Instancing generated Module: coreir.add(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__out;
  coreir_add #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$const_1_1__out;
  coreir_const #(.value(1'h1),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$const_1_1(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$const_1_1__out)
  );

  // Instancing generated Module: coreir.eq(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__out;
  coreir_eq #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1__out;
  coreir_const #(.value(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$const_1_1__out;
  coreir_const #(.value(1'h1),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$const_1_1(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$const_1_1__out)
  );

  // Instancing generated Module: coreir.add(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__out;
  coreir_add #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$const_1_1__out;
  coreir_const #(.value(1'h1),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$const_1_1(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$const_1_1__out)
  );

  // Instancing generated Module: coreir.eq(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__out;
  coreir_eq #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__in0;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__in1;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__sel;
  coreir_mux #(.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.const(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$const_0_2__out;
  coreir_const #(.value(2'h0),.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$const_0_2(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$const_0_2__out)
  );

  // Instancing generated Module: coreir.mux(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__in0;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__in1;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__sel;
  coreir_mux #(.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:2)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__clk;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__in;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out;
  coreir_reg #(.clk_posedge(1),.init(2'h0),.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out)
  );

  // Instancing generated Module: coreir.const(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$const_1_2__out;
  coreir_const #(.value(2'h1),.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$const_1_2(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$const_1_2__out)
  );

  // Instancing generated Module: coreir.add(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__in0;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__in1;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__out;
  coreir_add #(.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$const_2_2__out;
  coreir_const #(.value(2'h2),.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$const_2_2(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$const_2_2__out)
  );

  // Instancing generated Module: coreir.eq(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__in0;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__out;
  coreir_eq #(.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_const22_inst0__out;
  coreir_const #(.value(2'h2),.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_const22_inst0(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_const22_inst0__out)
  );

  // Instancing generated Module: coreir.eq(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__in0;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__out;
  coreir_eq #(.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__out)
  );

  // Instancing generated Module: coreir.ult(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__in0;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__out;
  coreir_ult #(.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__out)
  );

  // Instancing generated Module: coreir.mem(depth:2, has_init:False, width:8)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__raddr;
  wire [7:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__waddr;
  wire [7:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wen;
  coreir_mem #(.depth(2),.has_init(0),.width(8)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__clk),
    .raddr(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__raddr),
    .rdata(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata),
    .waddr(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__waddr),
    .wdata(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata),
    .wen(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wen)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1__out;
  coreir_const #(.value(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$const_1_1__out;
  coreir_const #(.value(1'h1),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$const_1_1(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$const_1_1__out)
  );

  // Instancing generated Module: coreir.add(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__out;
  coreir_add #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$const_1_1__out;
  coreir_const #(.value(1'h1),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$const_1_1(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$const_1_1__out)
  );

  // Instancing generated Module: coreir.eq(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__out;
  coreir_eq #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1__out;
  coreir_const #(.value(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$const_1_1__out;
  coreir_const #(.value(1'h1),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$const_1_1(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$const_1_1__out)
  );

  // Instancing generated Module: coreir.add(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__out;
  coreir_add #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$const_1_1__out;
  coreir_const #(.value(1'h1),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$const_1_1(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$const_1_1__out)
  );

  // Instancing generated Module: coreir.eq(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__out;
  coreir_eq #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__in0;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__in1;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__sel;
  coreir_mux #(.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.const(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$const_0_2__out;
  coreir_const #(.value(2'h0),.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$const_0_2(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$const_0_2__out)
  );

  // Instancing generated Module: coreir.mux(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__in0;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__in1;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__sel;
  coreir_mux #(.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:2)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__clk;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__in;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out;
  coreir_reg #(.clk_posedge(1),.init(2'h0),.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out)
  );

  // Instancing generated Module: coreir.const(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$const_1_2__out;
  coreir_const #(.value(2'h1),.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$const_1_2(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$const_1_2__out)
  );

  // Instancing generated Module: coreir.add(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__in0;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__in1;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__out;
  coreir_add #(.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$const_2_2__out;
  coreir_const #(.value(2'h2),.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$const_2_2(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$const_2_2__out)
  );

  // Instancing generated Module: coreir.eq(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__in0;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__out;
  coreir_eq #(.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_const22_inst0__out;
  coreir_const #(.value(2'h2),.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_const22_inst0(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_const22_inst0__out)
  );

  // Instancing generated Module: coreir.eq(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__in0;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__out;
  coreir_eq #(.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__out)
  );

  // Instancing generated Module: coreir.ult(width:2)
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__in0;
  wire [1:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__out;
  coreir_ult #(.width(2)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__out)
  );

  // Instancing generated Module: coreir.mem(depth:2, has_init:False, width:8)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__raddr;
  wire [7:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__waddr;
  wire [7:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wen;
  coreir_mem #(.depth(2),.has_init(0),.width(8)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__clk),
    .raddr(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__raddr),
    .rdata(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata),
    .waddr(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__waddr),
    .wdata(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata),
    .wen(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wen)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel;
  coreir_mux #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out),
    .sel(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0(
    .clk(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk),
    .in(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst0__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst0__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst1__in0;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst1__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst1__out;
  corebit_and TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst1(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst1__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst1__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst1__out)
  );

  // Instancing generated Module: coreir.const(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_const11_inst0__out;
  coreir_const #(.value(1'h1),.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_const11_inst0(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_const11_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:3)
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_const36_inst0__out;
  coreir_const #(.value(3'h6),.width(3)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_const36_inst0(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_const36_inst0__out)
  );

  // Instancing generated Module: coreir.eq(width:1)
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_1_inst0__in0;
  wire [0:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_1_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_1_inst0__out;
  coreir_eq #(.width(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_1_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_1_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_1_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_1_inst0__out)
  );

  // Instancing generated Module: coreir.eq(width:3)
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_3_inst0__in0;
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_3_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_3_inst0__out;
  coreir_eq #(.width(3)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_3_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_3_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_3_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_3_inst0__out)
  );

  // Instancing generated Module: coreir.ult(width:3)
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_ult3_inst0__in0;
  wire [2:0] TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_ult3_inst0__in1;
  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_ult3_inst0__out;
  coreir_ult #(.width(3)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_ult3_inst0(
    .in0(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_ult3_inst0__in0),
    .in1(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_ult3_inst0__in1),
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_ult3_inst0__out)
  );

  wire  TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$bit_const_1_None__out;
  corebit_const #(.value(1)) TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$bit_const_1_None(
    .out(TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$bit_const_1_None__out)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  wire  and_inst1__in0;
  wire  and_inst1__in1;
  wire  and_inst1__out;
  corebit_and and_inst1(
    .in0(and_inst1__in0),
    .in1(and_inst1__in1),
    .out(and_inst1__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] coreir_const81_inst0__out;
  coreir_const #(.value(8'h01),.width(8)) coreir_const81_inst0(
    .out(coreir_const81_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] coreir_const81_inst1__out;
  coreir_const #(.value(8'h01),.width(8)) coreir_const81_inst1(
    .out(coreir_const81_inst1__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] coreir_const81_inst2__out;
  coreir_const #(.value(8'h01),.width(8)) coreir_const81_inst2(
    .out(coreir_const81_inst2__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] coreir_const81_inst3__out;
  coreir_const #(.value(8'h01),.width(8)) coreir_const81_inst3(
    .out(coreir_const81_inst3__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] coreir_const82_inst0__out;
  coreir_const #(.value(8'h02),.width(8)) coreir_const82_inst0(
    .out(coreir_const82_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] coreir_const82_inst1__out;
  coreir_const #(.value(8'h02),.width(8)) coreir_const82_inst1(
    .out(coreir_const82_inst1__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] coreir_const82_inst2__out;
  coreir_const #(.value(8'h02),.width(8)) coreir_const82_inst2(
    .out(coreir_const82_inst2__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] coreir_const82_inst3__out;
  coreir_const #(.value(8'h02),.width(8)) coreir_const82_inst3(
    .out(coreir_const82_inst3__out)
  );

  // Instancing generated Module: coreir.mul(width:8)
  wire [7:0] coreir_mul8_inst0__in0;
  wire [7:0] coreir_mul8_inst0__in1;
  wire [7:0] coreir_mul8_inst0__out;
  coreir_mul #(.width(8)) coreir_mul8_inst0(
    .in0(coreir_mul8_inst0__in0),
    .in1(coreir_mul8_inst0__in1),
    .out(coreir_mul8_inst0__out)
  );

  // Instancing generated Module: coreir.mul(width:8)
  wire [7:0] coreir_mul8_inst1__in0;
  wire [7:0] coreir_mul8_inst1__in1;
  wire [7:0] coreir_mul8_inst1__out;
  coreir_mul #(.width(8)) coreir_mul8_inst1(
    .in0(coreir_mul8_inst1__in0),
    .in1(coreir_mul8_inst1__in1),
    .out(coreir_mul8_inst1__out)
  );

  // Instancing generated Module: coreir.mul(width:8)
  wire [7:0] coreir_mul8_inst2__in0;
  wire [7:0] coreir_mul8_inst2__in1;
  wire [7:0] coreir_mul8_inst2__out;
  coreir_mul #(.width(8)) coreir_mul8_inst2(
    .in0(coreir_mul8_inst2__in0),
    .in1(coreir_mul8_inst2__in1),
    .out(coreir_mul8_inst2__out)
  );

  // Instancing generated Module: coreir.mul(width:8)
  wire [7:0] coreir_mul8_inst3__in0;
  wire [7:0] coreir_mul8_inst3__in1;
  wire [7:0] coreir_mul8_inst3__out;
  coreir_mul #(.width(8)) coreir_mul8_inst3(
    .in0(coreir_mul8_inst3__in0),
    .in1(coreir_mul8_inst3__in1),
    .out(coreir_mul8_inst3__out)
  );

  // Instancing generated Module: coreir.mul(width:8)
  wire [7:0] coreir_mul8_inst4__in0;
  wire [7:0] coreir_mul8_inst4__in1;
  wire [7:0] coreir_mul8_inst4__out;
  coreir_mul #(.width(8)) coreir_mul8_inst4(
    .in0(coreir_mul8_inst4__in0),
    .in1(coreir_mul8_inst4__in1),
    .out(coreir_mul8_inst4__out)
  );

  // Instancing generated Module: coreir.mul(width:8)
  wire [7:0] coreir_mul8_inst5__in0;
  wire [7:0] coreir_mul8_inst5__in1;
  wire [7:0] coreir_mul8_inst5__out;
  coreir_mul #(.width(8)) coreir_mul8_inst5(
    .in0(coreir_mul8_inst5__in0),
    .in1(coreir_mul8_inst5__in1),
    .out(coreir_mul8_inst5__out)
  );

  // Instancing generated Module: coreir.mul(width:8)
  wire [7:0] coreir_mul8_inst6__in0;
  wire [7:0] coreir_mul8_inst6__in1;
  wire [7:0] coreir_mul8_inst6__out;
  coreir_mul #(.width(8)) coreir_mul8_inst6(
    .in0(coreir_mul8_inst6__in0),
    .in1(coreir_mul8_inst6__in1),
    .out(coreir_mul8_inst6__out)
  );

  // Instancing generated Module: coreir.mul(width:8)
  wire [7:0] coreir_mul8_inst7__in0;
  wire [7:0] coreir_mul8_inst7__in1;
  wire [7:0] coreir_mul8_inst7__out;
  coreir_mul #(.width(8)) coreir_mul8_inst7(
    .in0(coreir_mul8_inst7__in0),
    .in1(coreir_mul8_inst7__in1),
    .out(coreir_mul8_inst7__out)
  );

  assign ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_0_0$coreir_add8_inst0__in0[7:0] = ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_0$coreir_add8_inst0__out[7:0];

  assign ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_0_0$coreir_add8_inst0__in1[7:0] = ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_1$coreir_add8_inst0__out[7:0];

  assign O0[7:0] = ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_0_0$coreir_add8_inst0__out[7:0];

  assign ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_0$coreir_add8_inst0__in0[7:0] = coreir_mul8_inst0__out[7:0];

  assign ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_0$coreir_add8_inst0__in1[7:0] = coreir_mul8_inst1__out[7:0];

  assign ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_1$coreir_add8_inst0__in0[7:0] = coreir_mul8_inst2__out[7:0];

  assign ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst0$reducer$op_1_1$coreir_add8_inst0__in1[7:0] = coreir_mul8_inst3__out[7:0];

  assign ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_0_0$coreir_add8_inst0__in0[7:0] = ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_0$coreir_add8_inst0__out[7:0];

  assign ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_0_0$coreir_add8_inst0__in1[7:0] = ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_1$coreir_add8_inst0__out[7:0];

  assign O1[7:0] = ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_0_0$coreir_add8_inst0__out[7:0];

  assign ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_0$coreir_add8_inst0__in0[7:0] = coreir_mul8_inst4__out[7:0];

  assign ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_0$coreir_add8_inst0__in1[7:0] = coreir_mul8_inst5__out[7:0];

  assign ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_1$coreir_add8_inst0__in0[7:0] = coreir_mul8_inst6__out[7:0];

  assign ReduceParallel_n4_oprenamedForReduce_opcoreir_add8_I0_In_Bits_8___I1_In_Bits_8___O_Out_Bits_8____in0_In_Bits_8___in1_In_Bits_8___out_Out_Bits_8____inst1$reducer$op_1_1$coreir_add8_inst0__in1[7:0] = coreir_mul8_inst7__out[7:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join__in0[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$coreir_add3_inst0__out[2:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join__in1[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$const_0_3__out[2:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join__in1[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join__out[2:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$Mux2xOutBits3_inst0$coreir_commonlib_mux2x3_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join__in0[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__out[2:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__in[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join__out[2:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$enable_mux$coreir_commonlib_mux2x3_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$coreir_add3_inst0__in0[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__out[2:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$coreir_eq_3_inst0__in0[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__out[2:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_3_inst0__in0[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__out[2:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_ult3_inst0__in0[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_3_inst0$value__out[2:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$coreir_add3_inst0__in1[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$Counter3CER_inst0$const_1_3__out[2:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$and_inst0__in0 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$coreir_eq_3_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$and_inst0__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$coreir_eq_3_inst0__in1[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$Counter3_Mod7CE_inst0$const_6_3__out[2:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__in[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__waddr[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$const_1_1__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__in0 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$const_1_1__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__in[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__raddr[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$const_1_1__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__in0 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$const_1_1__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__in0[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__in1[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$const_0_2__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__in1[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__in0[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__in[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__in0[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__in0[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__in0[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__in0[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__in1[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$const_1_2__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__in0 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__in1[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$const_2_2__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__in0 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__in1[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_const22_inst0__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__in1[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_const22_inst0__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[1];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[2];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[3];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[4];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[5];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[6];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[7];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[1] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[2] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[3] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[4] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[5] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[6] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[7] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wen = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__in0 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__in1 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__in0 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__in1 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__in0 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I1[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst3__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst6__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I1[1];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst3__in0[1] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst6__in0[1] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I1[2];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst3__in0[2] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst6__in0[2] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I1[3];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst3__in0[3] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst6__in0[3] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I1[4];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst3__in0[4] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst6__in0[4] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I1[5];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst3__in0[5] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst6__in0[5] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I1[6];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst3__in0[6] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst6__in0[6] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I1[7];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst3__in0[7] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst6__in0[7] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst1__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst4__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst1__in0[1] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst4__in0[1] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst1__in0[2] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst4__in0[2] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst1__in0[3] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst4__in0[3] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst1__in0[4] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst4__in0[4] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst1__in0[5] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst4__in0[5] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst1__in0[6] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst4__in0[6] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst1__in0[7] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign coreir_mul8_inst4__in0[7] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst0$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__in[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__waddr[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$coreir_add1_inst0__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$Counter1CER_inst0$const_1_1__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__in0 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$and_inst0__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$coreir_eq_1_inst0__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst0$const_1_1__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$const_0_1__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$Mux2xOutBits1_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__in[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$enable_mux$coreir_commonlib_mux2x1_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__raddr[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0$value__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$coreir_add1_inst0__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$Counter1CER_inst0$const_1_1__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__in0 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$and_inst0__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$coreir_eq_1_inst0__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$Counter1_Mod2CE_inst1$const_1_1__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__in0[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__in1[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$const_0_2__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__in1[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$Mux2xOutBits2_inst0$coreir_commonlib_mux2x2_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__in0[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__in[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$enable_mux$coreir_commonlib_mux2x2_inst0$_join__sel = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__in0[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__in0[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__in0[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__in0[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_2_inst0$value__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$coreir_add2_inst0__in1[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$Counter2CER_inst0$const_1_2__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__in0 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$and_inst0__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$coreir_eq_2_inst0__in1[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$Counter2_Mod3CE_inst0$const_2_2__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__in0 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$and_inst0__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__in1[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_const22_inst0__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_ult2_inst0__in1[1:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_const22_inst0__out[1:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$InitialDelayCounter_2_inst0$coreir_eq_2_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[1];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[2];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[3];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[4];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[5];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[6];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__rdata[7];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[1] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[2] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[3] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[4] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[5] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[6] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wdata[7] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$NativeMapParallel_n1_opRAM_Array_8_In_Bit__t_2n_RADDR_In_Bits_1___RDATA_Array_8_Out_Bit___WADDR_In_Bits_1___WDATA_Array_8_In_Bit___WE_In_Bit__CLK_In_Clock___inst0$RAM_Array_8_In_Bit__t_2n_inst0$RAM2x8_inst0$coreir_mem2x8_inst0__wen = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__in0 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst0__in1 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__in0 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst1__in1 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$DelayedBuffer_Array_8_In_Bit__t_2n_1k_2emittingPeriod_2initialDelay_inst0$and_inst2__in0 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I0[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst7__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst2__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I0[1];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst7__in0[1] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst2__in0[1] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I0[2];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst7__in0[2] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst2__in0[2] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I0[3];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst7__in0[3] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst2__in0[3] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I0[4];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst7__in0[4] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst2__in0[4] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I0[5];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst7__in0[5] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst2__in0[5] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I0[6];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst7__in0[6] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst2__in0[6] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = I0[7];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst7__in0[7] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst2__in0[7] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_False_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst5__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst0__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_0$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst5__in0[1] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst0__in0[1] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_1$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst5__in0[2] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst0__in0[2] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_2$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst5__in0[3] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst0__in0[3] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_3$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst5__in0[4] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst0__in0[4] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_4$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst5__in0[5] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst0__in0[5] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_5$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst5__in0[6] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst0__in0[6] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_6$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__clk = CLK;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in1[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign coreir_mul8_inst5__in0[7] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst0$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__in0[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__in[0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$Mux2xNone_inst0$coreir_commonlib_mux2x1_inst0$_join__sel = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__clk = CLK;

  assign coreir_mul8_inst0__in0[7] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$NativeMapParallel_n1_opNativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___I_Array_2_Array_8_In_Bit____O_Array_2_Array_2_Array_2_Array_8_Out_Bit______CLK_Array_2_In_Clock___CE_Array_2_In_Enable____inst0$NativeMapParallel_n2_opshift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_I_Array_8_In_Bit___O_Array_2_Array_2_Array_8_Out_Bit_____CLK_In_Clock__CE_In_Enable___inst0$shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_inst1$shift_registers_for_shift_registers_for_AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_with__1_2__pxPerClock__8_8__imgSizes__2_2__neededCoordinates_True_lastInDimension_with__2__pxPerClock__8__imgSizes__2__neededCoordinates_True_lastInDimension_inst0$SIPO_Array_8_In_Bit__t_2n_0init_TrueCE_RESET_inst0$MapParallel_n8_opSIPO2CE_I_In_Bit__O_Out_Bits_2___CLK_In_Clock__CE_In_Enable___inst0$op_7$DFF_init0_has_ceTrue_has_resetFalse_has_async_resetFalse_inst1$reg_P_inst0__out[0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst0__in0 = and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst0__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_ult3_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst1__in0 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_1_inst0__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst1__in1 = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_3_inst0__out;

  assign valid_data_out = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$and_inst1__out;

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_1_inst0__in0[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_const11_inst0__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_1_inst0__in1[0:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_const11_inst0__out[0:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_eq_3_inst0__in1[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_const36_inst0__out[2:0];

  assign TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_ult3_inst0__in1[2:0] = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$AnyDimensionalLineBuffer_Array_8_In_Bit__type__1_2_pxPerClock__2_2_window__8_8_img__1_1_stride__0_0_origin_inst0$coreir_const36_inst0__out[2:0];

  assign ready_data_in = TwoDimensionalLineBuffer_Array_8_In_Bit__type_2x1pxPerClock_2x2window_8x8img_1x1stride_0x0origin_inst0$bit_const_1_None__out;

  assign and_inst0__in0 = valid_data_in;

  assign and_inst0__in1 = ready_data_out;

  assign and_inst1__in0 = and_inst0__out;

  assign and_inst1__in1 = CE;

  assign coreir_mul8_inst0__in1[7:0] = coreir_const81_inst0__out[7:0];

  assign coreir_mul8_inst4__in1[7:0] = coreir_const81_inst1__out[7:0];

  assign coreir_mul8_inst3__in1[7:0] = coreir_const81_inst2__out[7:0];

  assign coreir_mul8_inst7__in1[7:0] = coreir_const81_inst3__out[7:0];

  assign coreir_mul8_inst1__in1[7:0] = coreir_const82_inst0__out[7:0];

  assign coreir_mul8_inst5__in1[7:0] = coreir_const82_inst1__out[7:0];

  assign coreir_mul8_inst2__in1[7:0] = coreir_const82_inst2__out[7:0];

  assign coreir_mul8_inst6__in1[7:0] = coreir_const82_inst3__out[7:0];


endmodule  // partialParallel2Convolution_Circuit

